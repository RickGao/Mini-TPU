`default_nettype none
`timescale 1ns/1ns

module tpu (
    input wire clk,
    input wire rst_n,

    input wire [15:0] instruction,
    output wire [7:0] result
);



endmodule
